// DRV10975 Defines
`ifndef DRV10975_DEFINES
`define DRV10975_DEFINES

  `define SPEEDCTRL1    8'h00
  `define SPEEDCTRL2    8'h01
  `define DEVCTRL       8'h02
  `define EECTRL        8'h03
  `define STATUS        8'h10
  `define MOTORSPEED1   8'h11
  `define MOTORSPEED2   8'h12
  `define MOTORPERIOD1  8'h13
  `define MOTORPERIOD2  8'h14
  `define MOTORKT1      8'h15
  `define MOTORKT2      8'h16
  `define MOTORCURRENT1 8'h17
  `define MOTORCURRENT2 8'h18
  `define IPDPOSITION   8'h19
  `define SUPPLYVOLTAGE 8'h1A
  `define SPEEDCMD      8'h1B
  `define SPDCMDBUFFER  8'h1C
  `define FAULTCODE     8'h1E
  `define MOTORPARAM1   8'h20
  `define MOTORPARAM2   8'h21
  `define MOTORPARAM3   8'h22
  `define SYSOPT1       8'h23
  `define SYSOPT2       8'h24
  `define SYSOPT3       8'h25
  `define SYSOPT4       8'h26
  `define SYSOPT5       8'h27
  `define SYSOPT6       8'h28
  `define SYSOPT7       8'h29
  `define SYSOPT8       8'h2A
  `define SYSOPT9       8'h2B

  `define MOTORPARAM1_DEFAULT   8'h4A
  `define MOTORPARAM2_DEFAULT   8'h4E
  `define MOTORPARAM3_DEFAULT   8'h2A
  `define SYSOPT1_DEFAULT       8'h00
  `define SYSOPT2_DEFAULT       8'h98
  `define SYSOPT3_DEFAULT       8'hE4
  `define SYSOPT4_DEFAULT       8'h7A
  `define SYSOPT5_DEFAULT       8'hF4
  `define SYSOPT6_DEFAULT       8'h69
  `define SYSOPT7_DEFAULT       8'hB8
  `define SYSOPT8_DEFAULT       8'hAD
  `define SYSOPT9_DEFAULT       8'h0C

`endif

