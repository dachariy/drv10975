interface phase_if;
  reg U;
  reg V;
  reg W;
  reg FG;
endinterface
